module ex15 (
	input logic a, b, c, d,
	output logic y1, y2, y3
);

	
	
endmodule